module vtikz